module main;
initial begin
  $display("Hello, World!");
  $finish;
end
endmodule

===========================================
Created by: MD. Naiem Islam Nahid
File Type: Verilog
Magic Number: 2377
Time: 2024-11-07T04:57:22.486704
Date: Thursday, 07 November 2024, 2024th century
Emoji: None
===========================================
