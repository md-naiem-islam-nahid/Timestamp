module main;
initial begin
  $display("Hello, World!");
  $finish;
end
endmodule

===========================================
Created by: MD. Naiem Islam Nahid
File Type: Verilog
Magic Number: 5791
Time: 2024-11-07T05:02:54.290243
Date: Thursday, 07 November 2024, 2024th century
Emoji: None
===========================================
