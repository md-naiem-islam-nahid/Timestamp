library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity HelloWorld is
end HelloWorld;
architecture Behavioral of HelloWorld is
begin
process
begin
    report "Hello, World!";
    wait;
end process;
end Behavioral;

===========================================
Created by: MD. Naiem Islam Nahid
File Type: VHDL
Magic Number: 7395
Time: 2024-11-07T04:57:23.163889
Date: Thursday, 07 November 2024, 2024th century
Emoji: None
===========================================
